magic
tech sky130A
magscale 1 2
timestamp 1679710619
<< error_p >>
rect -173 536 -89 562
rect -173 530 197 536
rect 257 530 365 600
rect -209 494 221 500
rect -356 -541 -257 -373
rect -188 -540 -111 -328
rect 11 -540 88 -332
rect -188 -541 -83 -540
rect -23 -541 88 -540
rect -188 -545 88 -541
rect -188 -562 257 -545
rect -188 -582 256 -562
rect -183 -604 -177 -582
rect -89 -604 -83 -582
rect -183 -610 -83 -604
rect -23 -604 -17 -582
rect 11 -586 256 -582
rect 81 -604 87 -586
rect -23 -610 87 -604
<< nwell >>
rect -257 530 -173 562
rect 197 530 257 600
rect -257 -541 257 530
rect -257 -582 -188 -541
rect -111 -545 257 -541
rect -111 -582 11 -545
rect -257 -586 11 -582
rect 88 -562 257 -545
rect 88 -586 161 -562
rect -257 -600 161 -586
<< pmos >>
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
<< pdiff >>
rect -221 488 -159 500
rect -221 -488 -209 488
rect -175 -488 -159 488
rect -221 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 221 500
rect 159 -488 175 488
rect 209 -488 221 488
rect 159 -500 221 -488
<< pdiffc >>
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
<< poly >>
rect -159 500 -129 526
rect -63 500 -33 530
rect 33 500 63 526
rect 129 500 159 530
rect -159 -530 -129 -500
rect -63 -530 -33 -500
rect 33 -530 63 -500
rect 129 -530 159 -500
rect -223 -550 167 -530
rect -223 -590 -163 -550
rect -103 -590 7 -550
rect 67 -590 167 -550
rect -223 -620 167 -590
<< polycont >>
rect -163 -590 -103 -550
rect 7 -590 67 -550
<< locali >>
rect -209 488 -175 504
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -504 209 -488
<< viali >>
rect -209 81 -175 471
rect -113 -471 -79 -81
rect -17 81 17 471
rect 79 -471 113 -81
rect 175 81 209 471
rect -183 -550 -83 -540
rect -183 -590 -163 -550
rect -163 -590 -103 -550
rect -103 -590 -83 -550
rect -183 -610 -83 -590
rect -23 -550 87 -540
rect -23 -590 7 -550
rect 7 -590 67 -550
rect 67 -590 87 -550
rect -23 -610 87 -590
<< metal1 >>
rect -215 480 -169 483
rect -23 480 23 483
rect 169 480 215 483
rect -215 471 217 480
rect -215 81 -209 471
rect -175 81 -17 471
rect 17 81 175 471
rect 209 81 217 471
rect -215 80 217 81
rect -215 69 -169 80
rect -23 69 23 80
rect 169 69 215 80
rect -119 -80 -73 -69
rect 73 -80 119 -69
rect -119 -81 119 -80
rect -119 -471 -113 -81
rect -79 -470 79 -81
rect -79 -471 -73 -470
rect -119 -483 -73 -471
rect 73 -471 79 -470
rect 113 -471 119 -81
rect 73 -483 119 -471
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
