magic
tech sky130A
magscale 1 2
timestamp 1679528999
<< error_p >>
rect -29 1881 29 1887
rect -29 1847 -17 1881
rect -29 1841 29 1847
rect -29 -1847 29 -1841
rect -29 -1881 -17 -1847
rect -29 -1887 29 -1881
<< nwell >>
rect -211 -2019 211 2019
<< pmos >>
rect -15 -1800 15 1800
<< pdiff >>
rect -73 1788 -15 1800
rect -73 -1788 -61 1788
rect -27 -1788 -15 1788
rect -73 -1800 -15 -1788
rect 15 1788 73 1800
rect 15 -1788 27 1788
rect 61 -1788 73 1788
rect 15 -1800 73 -1788
<< pdiffc >>
rect -61 -1788 -27 1788
rect 27 -1788 61 1788
<< nsubdiff >>
rect -175 1949 -79 1983
rect 79 1949 175 1983
rect -175 1887 -141 1949
rect 141 1887 175 1949
rect -175 -1949 -141 -1887
rect 141 -1949 175 -1887
rect -175 -1983 -79 -1949
rect 79 -1983 175 -1949
<< nsubdiffcont >>
rect -79 1949 79 1983
rect -175 -1887 -141 1887
rect 141 -1887 175 1887
rect -79 -1983 79 -1949
<< poly >>
rect -33 1881 33 1897
rect -33 1847 -17 1881
rect 17 1847 33 1881
rect -33 1831 33 1847
rect -15 1800 15 1831
rect -15 -1831 15 -1800
rect -33 -1847 33 -1831
rect -33 -1881 -17 -1847
rect 17 -1881 33 -1847
rect -33 -1897 33 -1881
<< polycont >>
rect -17 1847 17 1881
rect -17 -1881 17 -1847
<< locali >>
rect -175 1949 -79 1983
rect 79 1949 175 1983
rect -175 1887 -141 1949
rect 141 1887 175 1949
rect -33 1847 -17 1881
rect 17 1847 33 1881
rect -61 1788 -27 1804
rect -61 -1804 -27 -1788
rect 27 1788 61 1804
rect 27 -1804 61 -1788
rect -33 -1881 -17 -1847
rect 17 -1881 33 -1847
rect -175 -1949 -141 -1887
rect 141 -1949 175 -1887
rect -175 -1983 -79 -1949
rect 79 -1983 175 -1949
<< viali >>
rect -17 1847 17 1881
rect -61 -1788 -27 1788
rect 27 -1788 61 1788
rect -17 -1881 17 -1847
<< metal1 >>
rect -29 1881 29 1887
rect -29 1847 -17 1881
rect 17 1847 29 1881
rect -29 1841 29 1847
rect -67 1788 -21 1800
rect -67 -1788 -61 1788
rect -27 -1788 -21 1788
rect -67 -1800 -21 -1788
rect 21 1788 67 1800
rect 21 -1788 27 1788
rect 61 -1788 67 1788
rect 21 -1800 67 -1788
rect -29 -1847 29 -1841
rect -29 -1881 -17 -1847
rect 17 -1881 29 -1847
rect -29 -1887 29 -1881
<< properties >>
string FIXED_BBOX -158 -1966 158 1966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 18.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
