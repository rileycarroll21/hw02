magic
tech sky130A
magscale 1 2
timestamp 1679633613
<< error_p >>
rect -257 520 257 536
rect -221 484 221 500
<< nwell >>
rect -257 -584 257 520
<< pmos >>
rect -159 -500 -127 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
<< pdiff >>
rect -221 488 -159 500
rect -221 -488 -209 488
rect -175 -488 -159 488
rect -221 -500 -159 -488
rect -127 488 -63 500
rect -127 -488 -113 488
rect -79 -488 -63 488
rect -127 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 221 500
rect 159 -488 175 488
rect 209 -488 221 488
rect 159 -500 221 -488
<< pdiffc >>
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
<< poly >>
rect -159 500 -127 520
rect -63 500 -33 520
rect 33 500 63 520
rect 129 500 159 520
rect -159 -524 -127 -500
rect -63 -524 -33 -500
rect 33 -524 63 -500
rect 129 -524 159 -500
rect -223 -554 217 -524
rect -223 -604 -173 -554
rect -113 -604 -23 -554
rect 37 -604 117 -554
rect 177 -604 217 -554
rect -223 -624 217 -604
<< polycont >>
rect -173 -604 -113 -554
rect -23 -604 37 -554
rect 117 -604 177 -554
<< locali >>
rect -209 488 -175 504
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -504 209 -488
<< viali >>
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect -193 -554 -93 -544
rect -193 -604 -173 -554
rect -173 -604 -113 -554
rect -113 -604 -93 -554
rect -193 -614 -93 -604
rect -43 -554 57 -544
rect -43 -604 -23 -554
rect -23 -604 37 -554
rect 37 -604 57 -554
rect -43 -614 57 -604
rect 97 -554 197 -544
rect 97 -604 117 -554
rect 117 -604 177 -554
rect 177 -604 197 -554
rect 97 -614 197 -604
<< metal1 >>
rect -215 488 -169 500
rect -215 -488 -209 488
rect -175 -488 -169 488
rect -215 -500 -169 -488
rect -119 488 -73 500
rect -119 -488 -113 488
rect -79 -488 -73 488
rect -119 -500 -73 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 73 488 119 500
rect 73 -488 79 488
rect 113 -488 119 488
rect 73 -500 119 -488
rect 169 488 215 500
rect 169 -488 175 488
rect 209 -488 215 488
rect 169 -500 215 -488
rect -223 -544 217 -534
rect -223 -614 -193 -544
rect -93 -614 -43 -544
rect 57 -614 97 -544
rect 197 -614 217 -544
rect -223 -624 217 -614
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
