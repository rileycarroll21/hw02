magic
tech sky130A
timestamp 1679555532
<< error_p >>
rect -18 286 18 289
rect -18 269 -12 286
rect -18 266 18 269
rect -18 -269 18 -266
rect -18 -286 -12 -269
rect -18 -289 18 -286
<< pwell >>
rect -118 -355 118 355
<< nmos >>
rect -20 -250 20 250
<< ndiff >>
rect -49 244 -20 250
rect -49 -244 -43 244
rect -26 -244 -20 244
rect -49 -250 -20 -244
rect 20 244 49 250
rect 20 -244 26 244
rect 43 -244 49 244
rect 20 -250 49 -244
<< ndiffc >>
rect -43 -244 -26 244
rect 26 -244 43 244
<< psubdiff >>
rect -100 320 -52 337
rect 52 320 100 337
rect -100 289 -83 320
rect 83 289 100 320
rect -100 -320 -83 -289
rect 83 -320 100 -289
rect -100 -337 -52 -320
rect 52 -337 100 -320
<< psubdiffcont >>
rect -52 320 52 337
rect -100 -289 -83 289
rect 83 -289 100 289
rect -52 -337 52 -320
<< poly >>
rect -20 286 20 294
rect -20 269 -12 286
rect 12 269 20 286
rect -20 250 20 269
rect -20 -269 20 -250
rect -20 -286 -12 -269
rect 12 -286 20 -269
rect -20 -294 20 -286
<< polycont >>
rect -12 269 12 286
rect -12 -286 12 -269
<< locali >>
rect -100 320 -52 337
rect 52 320 100 337
rect -100 289 -83 320
rect 83 289 100 320
rect -20 269 -12 286
rect 12 269 20 286
rect -43 244 -26 252
rect -43 -252 -26 -244
rect 26 244 43 252
rect 26 -252 43 -244
rect -20 -286 -12 -269
rect 12 -286 20 -269
rect -100 -320 -83 -289
rect 83 -320 100 -289
rect -100 -337 -52 -320
rect 52 -337 100 -320
<< viali >>
rect -12 269 12 286
rect -43 -244 -26 244
rect 26 -244 43 244
rect -12 -286 12 -269
<< metal1 >>
rect -18 286 18 289
rect -18 269 -12 286
rect 12 269 18 286
rect -18 266 18 269
rect -46 244 -23 250
rect -46 -244 -43 244
rect -26 -244 -23 244
rect -46 -250 -23 -244
rect 23 244 46 250
rect 23 -244 26 244
rect 43 -244 46 244
rect 23 -250 46 -244
rect -18 -269 18 -266
rect -18 -286 -12 -269
rect 12 -286 18 -269
rect -18 -289 18 -286
<< properties >>
string FIXED_BBOX -91 -328 91 328
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
