magic
tech sky130A
magscale 1 2
timestamp 1679530569
<< error_p >>
rect 6280 2453 6338 2459
rect 6326 2419 6338 2453
rect 6280 2413 6338 2419
<< error_s >>
rect -2387 6126 -2341 6138
rect 1741 6126 1787 6138
rect -2387 6092 -2381 6126
rect 1741 6092 1747 6126
rect -2387 6080 -2341 6092
rect 1741 6080 1787 6092
rect 1900 6000 2054 6218
rect 5946 6200 6100 6218
rect 6041 6126 6087 6138
rect 6041 6092 6047 6126
rect 6041 6080 6087 6092
rect 6200 6000 6354 6200
rect -2390 5690 -2344 5702
rect 1720 5690 1766 5702
rect 1910 5690 1956 5702
rect 6020 5690 6066 5702
rect -2390 5656 -2384 5690
rect 1720 5656 1726 5690
rect 1910 5656 1916 5690
rect 6020 5656 6026 5690
rect -2390 5644 -2344 5656
rect 1720 5644 1766 5656
rect 1910 5644 1956 5656
rect 6020 5644 6066 5656
rect -390 4322 -344 4334
rect 720 4322 766 4334
rect -390 4274 -384 4322
rect 720 4274 726 4322
rect -390 4262 -344 4274
rect 720 4262 766 4274
use sky130_fd_pr__nfet_01v8_P64V6L  XM1
timestamp 1679529196
transform 0 -1 -1812 1 0 4363
box -163 -588 163 588
use sky130_fd_pr__nfet_01v8_QREW3P  XM2
timestamp 1679529196
transform 0 -1 188 1 0 4298
box -98 -588 98 588
use sky130_fd_pr__pfet_01v8_MGSX2X  XM3
timestamp 1679530569
transform 0 -1 -300 1 0 6109
box -109 -2100 109 2100
use sky130_fd_pr__nfet_01v8_YMW3AY  XM5
timestamp 1679529196
transform 0 -1 -312 1 0 5673
box -73 -2088 73 2088
use sky130_fd_pr__pfet_01v8_XGSKWQ  XM7
timestamp 1679529196
transform -1 0 6309 0 -1 4300
box -109 -1900 109 1900
use sky130_fd_pr__nfet_01v8_VB4QDD  XM8
timestamp 1679529196
transform 0 -1 1563 1 0 4333
box -133 -163 133 163
use sky130_fd_pr__nfet_01v8_YMW3AY  sky130_fd_pr__nfet_01v8_YMW3AY_0
timestamp 1679529196
transform 0 -1 3988 1 0 5673
box -73 -2088 73 2088
use sky130_fd_pr__pfet_01v8_MGSX2X  sky130_fd_pr__pfet_01v8_MGSX2X_0
timestamp 1679530569
transform 0 -1 4000 1 0 6109
box -109 -2100 109 2100
<< end >>
