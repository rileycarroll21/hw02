magic
tech sky130A
magscale 1 2
timestamp 1679889462
<< nwell >>
rect -1100 3900 3000 5200
<< psubdiff >>
rect 2116 3180 2140 3420
rect 2680 3180 2704 3420
rect -2244 1740 -2220 2320
rect 220 1740 244 2320
<< nsubdiff >>
rect -160 5000 880 5060
rect -160 4700 -100 5000
rect 800 4700 880 5000
rect -160 4660 880 4700
rect 1300 5020 2340 5060
rect 1300 4680 1340 5020
rect 2300 4680 2340 5020
rect 1300 4660 2340 4680
<< psubdiffcont >>
rect 2140 3180 2680 3420
rect -2220 1740 220 2320
<< nsubdiffcont >>
rect -100 4700 800 5000
rect 1340 4680 2300 5020
<< locali >>
rect -660 5060 2800 5100
rect -660 4660 -160 5060
rect 880 5020 2800 5060
rect 880 4660 1320 5020
rect 2320 4660 2800 5020
rect -660 4600 2800 4660
rect 2340 3437 2460 3540
rect 2124 3180 2131 3420
rect -2140 2320 -1180 2540
rect -820 2320 140 2600
rect -2236 1740 -2220 2320
rect 220 1740 236 2320
<< viali >>
rect -160 5000 880 5060
rect -160 4700 -100 5000
rect -100 4700 800 5000
rect 800 4700 880 5000
rect -160 4660 880 4700
rect 1320 4680 1340 5020
rect 1340 4680 2300 5020
rect 2300 4680 2320 5020
rect 1320 4660 2320 4680
rect 2131 3420 2702 3437
rect 2131 3180 2140 3420
rect 2140 3180 2680 3420
rect 2680 3180 2702 3420
rect 2131 3178 2702 3180
rect -2207 1746 167 2300
<< metal1 >>
rect -1820 5060 3340 5100
rect -1820 4660 -160 5060
rect 880 5020 3340 5060
rect 880 4660 1320 5020
rect 2320 4660 3340 5020
rect -1820 4620 3340 4660
rect -1820 3020 -1400 4620
rect -920 4430 -510 4620
rect -360 4050 40 4380
rect -250 3960 40 4050
rect 90 4040 520 4470
rect 580 4130 950 4620
rect 137 4035 517 4040
rect 200 3960 460 4035
rect -250 3720 460 3960
rect 1120 3960 1520 4180
rect 1620 4040 1880 4460
rect 1920 4400 2280 4620
rect 2340 4040 2680 4380
rect 1620 3960 1780 4040
rect 1120 3720 1780 3960
rect 2340 3740 2520 4040
rect -1040 3220 -870 3680
rect -250 3630 150 3720
rect -690 3500 -400 3580
rect -680 3100 -410 3500
rect 520 3100 900 3480
rect 1120 3360 1460 3720
rect 2960 3700 3340 4620
rect 1520 3240 1780 3680
rect 2520 3560 3340 3700
rect 2336 3450 2452 3538
rect 2101 3437 2711 3450
rect 2101 3400 2131 3437
rect -1820 2860 -860 3020
rect -1820 2800 -1400 2860
rect -1120 2600 -860 2860
rect -680 2840 900 3100
rect 2100 3178 2131 3400
rect 2702 3178 2711 3437
rect 2100 3061 2711 3178
rect -680 2720 140 2840
rect -2020 2331 -1330 2560
rect -630 2331 60 2610
rect -2233 2330 207 2331
rect 2100 2330 2700 3061
rect -2233 2300 2700 2330
rect -2233 1766 -2207 2300
rect -2237 1746 -2207 1766
rect 167 1750 2700 2300
rect 167 1746 255 1750
rect -2237 1720 255 1746
use sky130_fd_pr__nfet_01v8_P64V6L  XM1
timestamp 1679639255
transform 0 -1 -1659 1 0 2675
box -163 -588 163 528
use sky130_fd_pr__nfet_01v8_QREW3P  XM2
timestamp 1679638617
transform 0 -1 -328 1 0 2666
box -98 -532 102 608
use sky130_fd_pr__nfet_01v8_L7MCXF  XM5
timestamp 1679699828
transform 0 1 -332 -1 0 3461
box -239 -628 221 526
use sky130_fd_pr__pfet_01v8_FBJWLQ  XM7
timestamp 1679810962
transform 0 -1 2350 1 0 4257
box -355 -550 347 701
use sky130_fd_pr__nfet_01v8_8C4LHH  XM8
timestamp 1679640193
transform 0 1 2432 -1 0 3633
box -133 -132 133 132
use sky130_fd_pr__nfet_01v8_L7MCXF  sky130_fd_pr__nfet_01v8_L7MCXF_0
timestamp 1679699828
transform 0 -1 1006 1 0 3499
box -239 -628 221 526
use sky130_fd_pr__pfet_01v8_CQ5Q4H  sky130_fd_pr__pfet_01v8_CQ5Q4H_0
timestamp 1679710619
transform 0 1 1040 -1 0 4257
box -356 -620 365 600
use sky130_fd_pr__pfet_01v8_CQ5Q4H  sky130_fd_pr__pfet_01v8_CQ5Q4H_1
timestamp 1679710619
transform 0 -1 -437 1 0 4265
box -356 -620 365 600
<< labels >>
rlabel metal1 -1000 3280 -920 3620 1 in_p
port 6 n
rlabel locali -640 2410 -390 2510 1 Vss
port 8 n
rlabel metal1 2340 3780 2520 4000 1 amp_out
port 4 n
rlabel metal1 1540 3260 1740 3620 1 in_n
port 5 n
rlabel nwell -160 4660 880 5060 1 Vdd
port 7 n
<< end >>
