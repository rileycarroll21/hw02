magic
tech sky130A
magscale 1 2
timestamp 1679530569
<< error_p >>
rect -29 2081 29 2087
rect -29 2047 -17 2081
rect -29 2041 29 2047
rect -29 -2047 29 -2041
rect -29 -2081 -17 -2047
rect -29 -2087 29 -2081
<< nwell >>
rect -109 -2100 109 2100
<< pmos >>
rect -15 -2000 15 2000
<< pdiff >>
rect -73 1988 -15 2000
rect -73 -1988 -61 1988
rect -27 -1988 -15 1988
rect -73 -2000 -15 -1988
rect 15 1988 73 2000
rect 15 -1988 27 1988
rect 61 -1988 73 1988
rect 15 -2000 73 -1988
<< pdiffc >>
rect -61 -1988 -27 1988
rect 27 -1988 61 1988
<< poly >>
rect -33 2081 33 2097
rect -33 2047 -17 2081
rect 17 2047 33 2081
rect -33 2031 33 2047
rect -15 2000 15 2031
rect -15 -2031 15 -2000
rect -33 -2047 33 -2031
rect -33 -2081 -17 -2047
rect 17 -2081 33 -2047
rect -33 -2097 33 -2081
<< polycont >>
rect -17 2047 17 2081
rect -17 -2081 17 -2047
<< locali >>
rect -33 2047 -17 2081
rect 17 2047 33 2081
rect -61 1988 -27 2004
rect -61 -2004 -27 -1988
rect 27 1988 61 2004
rect 27 -2004 61 -1988
rect -33 -2081 -17 -2047
rect 17 -2081 33 -2047
<< viali >>
rect -17 2047 17 2081
rect -61 -1988 -27 1988
rect 27 -1988 61 1988
rect -17 -2081 17 -2047
<< metal1 >>
rect -29 2081 29 2087
rect -29 2047 -17 2081
rect 17 2047 29 2081
rect -29 2041 29 2047
rect -67 1988 -21 2000
rect -67 -1988 -61 1988
rect -27 -1988 -21 1988
rect -67 -2000 -21 -1988
rect 21 1988 67 2000
rect 21 -1988 27 1988
rect 61 -1988 67 1988
rect 21 -2000 67 -1988
rect -29 -2047 29 -2041
rect -29 -2081 -17 -2047
rect 17 -2081 29 -2047
rect -29 -2087 29 -2081
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
