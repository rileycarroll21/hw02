magic
tech sky130A
magscale 1 2
timestamp 1679555532
<< error_p >>
rect -77 531 -19 537
rect 115 531 173 537
rect -77 497 -65 531
rect 115 497 127 531
rect -77 491 -19 497
rect 115 491 173 497
rect -173 -497 -115 -491
rect 19 -497 77 -491
rect -173 -531 -161 -497
rect 19 -531 31 -497
rect -173 -537 -115 -531
rect 19 -537 77 -531
<< nwell >>
rect -359 -669 359 669
<< pmos >>
rect -159 -450 -129 450
rect -63 -450 -33 450
rect 33 -450 63 450
rect 129 -450 159 450
<< pdiff >>
rect -221 438 -159 450
rect -221 -438 -209 438
rect -175 -438 -159 438
rect -221 -450 -159 -438
rect -129 438 -63 450
rect -129 -438 -113 438
rect -79 -438 -63 438
rect -129 -450 -63 -438
rect -33 438 33 450
rect -33 -438 -17 438
rect 17 -438 33 438
rect -33 -450 33 -438
rect 63 438 129 450
rect 63 -438 79 438
rect 113 -438 129 438
rect 63 -450 129 -438
rect 159 438 221 450
rect 159 -438 175 438
rect 209 -438 221 438
rect 159 -450 221 -438
<< pdiffc >>
rect -209 -438 -175 438
rect -113 -438 -79 438
rect -17 -438 17 438
rect 79 -438 113 438
rect 175 -438 209 438
<< nsubdiff >>
rect -323 599 -227 633
rect 227 599 323 633
rect -323 537 -289 599
rect 289 537 323 599
rect -323 -599 -289 -537
rect 289 -599 323 -537
rect -323 -633 -227 -599
rect 227 -633 323 -599
<< nsubdiffcont >>
rect -227 599 227 633
rect -323 -537 -289 537
rect 289 -537 323 537
rect -227 -633 227 -599
<< poly >>
rect -81 531 -15 547
rect -81 497 -65 531
rect -31 497 -15 531
rect -81 481 -15 497
rect 111 531 177 547
rect 111 497 127 531
rect 161 497 177 531
rect 111 481 177 497
rect -159 450 -129 476
rect -63 450 -33 481
rect 33 450 63 476
rect 129 450 159 481
rect -159 -481 -129 -450
rect -63 -476 -33 -450
rect 33 -481 63 -450
rect 129 -476 159 -450
rect -177 -497 -111 -481
rect -177 -531 -161 -497
rect -127 -531 -111 -497
rect -177 -547 -111 -531
rect 15 -497 81 -481
rect 15 -531 31 -497
rect 65 -531 81 -497
rect 15 -547 81 -531
<< polycont >>
rect -65 497 -31 531
rect 127 497 161 531
rect -161 -531 -127 -497
rect 31 -531 65 -497
<< locali >>
rect -323 599 -227 633
rect 227 599 323 633
rect -323 537 -289 599
rect 289 537 323 599
rect -81 497 -65 531
rect -31 497 -15 531
rect 111 497 127 531
rect 161 497 177 531
rect -209 438 -175 454
rect -209 -454 -175 -438
rect -113 438 -79 454
rect -113 -454 -79 -438
rect -17 438 17 454
rect -17 -454 17 -438
rect 79 438 113 454
rect 79 -454 113 -438
rect 175 438 209 454
rect 175 -454 209 -438
rect -177 -531 -161 -497
rect -127 -531 -111 -497
rect 15 -531 31 -497
rect 65 -531 81 -497
rect -323 -599 -289 -537
rect 289 -599 323 -537
rect -323 -633 -227 -599
rect 227 -633 323 -599
<< viali >>
rect -65 497 -31 531
rect 127 497 161 531
rect -209 -438 -175 438
rect -113 -438 -79 438
rect -17 -438 17 438
rect 79 -438 113 438
rect 175 -438 209 438
rect -161 -531 -127 -497
rect 31 -531 65 -497
<< metal1 >>
rect -77 531 -19 537
rect -77 497 -65 531
rect -31 497 -19 531
rect -77 491 -19 497
rect 115 531 173 537
rect 115 497 127 531
rect 161 497 173 531
rect 115 491 173 497
rect -215 438 -169 450
rect -215 -438 -209 438
rect -175 -438 -169 438
rect -215 -450 -169 -438
rect -119 438 -73 450
rect -119 -438 -113 438
rect -79 -438 -73 438
rect -119 -450 -73 -438
rect -23 438 23 450
rect -23 -438 -17 438
rect 17 -438 23 438
rect -23 -450 23 -438
rect 73 438 119 450
rect 73 -438 79 438
rect 113 -438 119 438
rect 73 -450 119 -438
rect 169 438 215 450
rect 169 -438 175 438
rect 209 -438 215 438
rect 169 -450 215 -438
rect -173 -497 -115 -491
rect -173 -531 -161 -497
rect -127 -531 -115 -497
rect -173 -537 -115 -531
rect 19 -497 77 -491
rect 19 -531 31 -497
rect 65 -531 77 -497
rect 19 -537 77 -531
<< properties >>
string FIXED_BBOX -306 -616 306 616
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.5 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
