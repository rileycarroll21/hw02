magic
tech sky130A
magscale 1 2
timestamp 1679555532
<< error_p >>
rect -77 572 -19 578
rect 115 572 173 578
rect -77 538 -65 572
rect 115 538 127 572
rect -77 532 -19 538
rect 115 532 173 538
rect -173 -538 -115 -532
rect 19 -538 77 -532
rect -173 -572 -161 -538
rect 19 -572 31 -538
rect -173 -578 -115 -572
rect 19 -578 77 -572
<< pwell >>
rect -359 -710 359 710
<< nmos >>
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
<< ndiff >>
rect -221 488 -159 500
rect -221 -488 -209 488
rect -175 -488 -159 488
rect -221 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 221 500
rect 159 -488 175 488
rect 209 -488 221 488
rect 159 -500 221 -488
<< ndiffc >>
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
<< psubdiff >>
rect -323 640 -227 674
rect 227 640 323 674
rect -323 578 -289 640
rect 289 578 323 640
rect -323 -640 -289 -578
rect 289 -640 323 -578
rect -323 -674 -227 -640
rect 227 -674 323 -640
<< psubdiffcont >>
rect -227 640 227 674
rect -323 -578 -289 578
rect 289 -578 323 578
rect -227 -674 227 -640
<< poly >>
rect -81 572 -15 588
rect -81 538 -65 572
rect -31 538 -15 572
rect -159 500 -129 526
rect -81 522 -15 538
rect 111 572 177 588
rect 111 538 127 572
rect 161 538 177 572
rect -63 500 -33 522
rect 33 500 63 526
rect 111 522 177 538
rect 129 500 159 522
rect -159 -522 -129 -500
rect -177 -538 -111 -522
rect -63 -526 -33 -500
rect 33 -522 63 -500
rect -177 -572 -161 -538
rect -127 -572 -111 -538
rect -177 -588 -111 -572
rect 15 -538 81 -522
rect 129 -526 159 -500
rect 15 -572 31 -538
rect 65 -572 81 -538
rect 15 -588 81 -572
<< polycont >>
rect -65 538 -31 572
rect 127 538 161 572
rect -161 -572 -127 -538
rect 31 -572 65 -538
<< locali >>
rect -323 640 -227 674
rect 227 640 323 674
rect -323 578 -289 640
rect 289 578 323 640
rect -81 538 -65 572
rect -31 538 -15 572
rect 111 538 127 572
rect 161 538 177 572
rect -209 488 -175 504
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -504 209 -488
rect -177 -572 -161 -538
rect -127 -572 -111 -538
rect 15 -572 31 -538
rect 65 -572 81 -538
rect -323 -640 -289 -578
rect 289 -640 323 -578
rect -323 -674 -227 -640
rect 227 -674 323 -640
<< viali >>
rect -65 538 -31 572
rect 127 538 161 572
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect -161 -572 -127 -538
rect 31 -572 65 -538
<< metal1 >>
rect -77 572 -19 578
rect -77 538 -65 572
rect -31 538 -19 572
rect -77 532 -19 538
rect 115 572 173 578
rect 115 538 127 572
rect 161 538 173 572
rect 115 532 173 538
rect -215 488 -169 500
rect -215 -488 -209 488
rect -175 -488 -169 488
rect -215 -500 -169 -488
rect -119 488 -73 500
rect -119 -488 -113 488
rect -79 -488 -73 488
rect -119 -500 -73 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 73 488 119 500
rect 73 -488 79 488
rect 113 -488 119 488
rect 73 -500 119 -488
rect 169 488 215 500
rect 169 -488 175 488
rect 209 -488 215 488
rect 169 -500 215 -488
rect -173 -538 -115 -532
rect -173 -572 -161 -538
rect -127 -572 -115 -538
rect -173 -578 -115 -572
rect 19 -538 77 -532
rect 19 -572 31 -538
rect 65 -572 77 -538
rect 19 -578 77 -572
<< properties >>
string FIXED_BBOX -306 -657 306 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
